module lab4iram2F(CLK, RESET, ADDR, Q);
  input         CLK;
  input         RESET;
  input  [7:0]  ADDR;
  output [15:0] Q;

  reg    [15:0] mem[0:127]; // instruction memory with 16 bit entries

  wire   [6:0]  saddr;
  integer       i;

  assign saddr = ADDR[7:1];
  assign Q = mem[saddr];

  always @(posedge CLK) begin
    if(RESET) begin

      mem[0] <= 16'b1111000000000001; //   SUB R0, R0, R0
      mem[1] <= 16'b0000000000000001; //   HALT
      mem[2] <= 16'b1111010010010001; //   SUB R2, R2, R2
      mem[3] <= 16'b0000000000000000; //   ADDI R4, R2, -30
      mem[4] <= 16'b1011100000000001; //   BLTZ R4, 1
      mem[5] <= 16'b0101000010011101; //   ADDI R2, R0, 29
      mem[6] <= 16'b1111010000010100; //   SLL R2, R2
      mem[7] <= 16'b1111011011011001; //   SUB R3, R3, R3
      mem[8] <= 16'b0100000011111110; //   SB R3, -2(R0)
      mem[9] <= 16'b0010000011111001; //   LB R3, -2(R0)
      mem[10] <= 16'b0100000011111111; //   SB R3, -1(R0)
      mem[11] <= 16'b0101000001100000; //   ADDI R1, R0,-32
      mem[12] <= 16'b1111001000001100; //   SLL R1,R1
      mem[13] <= 16'b1111001000001100; //   SLL R1, R1
      mem[14] <= 16'b0101000101000110; //   ADDI R5, R0, 6
      mem[15] <= 16'b1111101010101001; //   SUB R5, R5, R2
      mem[16] <= 16'b1011101000010101; //   BLTZ R5, 21
      mem[17] <= 16'b0101000101000110; //   ADDI R5, R0, 6
      mem[18] <= 16'b1001010101010010; //   BNE R5, R2, 18
      mem[19] <= 16'b0110000101000111; //   ANDI R5, R0, 7
      mem[20] <= 16'b1111001000001010; //   SRA R1, R1
      mem[21] <= 16'b1000010101001111; //   BEQ R5, R2, 15
      mem[22] <= 16'b0101000101001000; //   ADDI R5, R0, 8
      mem[23] <= 16'b1111001000001010; //   SRA R1, R1
      mem[24] <= 16'b1000010101001100; //   BEQ R5, R2, 12
      mem[25] <= 16'b0101000101001001; //   ADDI R5, R0, 9
      mem[26] <= 16'b1111001000001010; //   SRA R1, R1
      mem[27] <= 16'b1001010101001001; //   BNE R5, R2, 9
      mem[28] <= 16'b0110000101001010; //   ANDI R5, R0, 10
      mem[29] <= 16'b1111001000001010; //   SRA R1, R1
      mem[30] <= 16'b1000010101000110; //   BEQ R5, R2, 6
      mem[31] <= 16'b0101000101001011; //   ADDI R5, R0, 11
      mem[32] <= 16'b1111001000001010; //   SRA R1, R1
      mem[33] <= 16'b1001010101000011; //   BNE R5, R2, 3
      mem[34] <= 16'b0101000101001100; //   ADDI R5, R0, 12
      mem[35] <= 16'b1111001000001010; //   SRA R1, R1
      mem[36] <= 16'b1000010101000001; //   BEQ R5, R2, 1
      mem[37] <= 16'b1111001000001010; //   SRA R1,R1
      mem[38] <= 16'b0100000001111100; //   SB R1, -4(R0)

      for(i = 39; i < 128; i = i + 1) begin
        mem[i] <= 16'b0000000000000000;
      end
    end
  end

endmodule