module lab4iramHRMmod(CLK, RESET, ADDR, Q);
  input         CLK;
  input         RESET;
  input  [7:0]  ADDR;
  output [15:0] Q;

  reg    [15:0] mem[0:127]; // instruction memory with 16 bit entries

  wire   [6:0]  saddr;
  integer       i;

  assign saddr = ADDR[7:1];
  assign Q = mem[saddr];

  always @(posedge CLK) begin
    if(RESET) begin

      // data goes here
      mem[0] <= 16'b1111000000000001; //   SUB R0, R0, R0
      mem[1] <= 16'b1111010010010001; //   SUB R2, R2, R2
      mem[2] <= 16'b1111111111111001; //   SUB R7, R7, R7
      mem[3] <= 16'b1111110110110001; //   SUB R6, R6, R6
      mem[4] <= 16'b0101000101111111; //   ADDI R5, R0, -1
      mem[5] <= 16'b1111101000101011; //   SRL R5, R5
      mem[6] <= 16'b0010000011111011; //   LB R3, -5(R0)
      mem[7] <= 16'b0110011011000001; //   ANDI R3, R3, 1
      mem[8] <= 16'b0010000100111011; //   LB R4, -5(R0)
      mem[9] <= 16'b0110100100000001; //   ANDI R4, R4, 1
      mem[10] <= 16'b1111100011011000; //   ADD R3, R4, R3
      mem[11] <= 16'b0110011011000001; //   ANDI R3, R3, 1
      mem[12] <= 16'b1111011100011101; //   AND R3, R3, R4
      mem[13] <= 16'b1111010011010000; //   ADD R2, R2, R3
      mem[14] <= 16'b1111100000011000; //   ADD R3, R4, R0
      mem[15] <= 16'b0101111111111111; //   ADDI R7, R7, -1
      mem[16] <= 16'b1001000111110111; //   BNE R7, R0, -9
      mem[17] <= 16'b0101110110111111; //   ADDI R6, R6, -1
      mem[18] <= 16'b1001000110110101; //   BNE R6, R0, -11
      mem[19] <= 16'b0101101101111111; //   ADDI R5, R5, -1
      mem[20] <= 16'b1001000101110011; //   BNE R5, R0, -13
      mem[21] <= 16'b0101010100100010; //   ADDI R4, R2, -30
      mem[22] <= 16'b1011100000000001; //   BLTZ R4, 1
      mem[23] <= 16'b0101000010011101; //   ADDI R2, R0, 29
      mem[24] <= 16'b1111010000010100; //   SLL R2, R2
      mem[25] <= 16'b0010010011000000; //   LB R3, 0(R2)
      mem[26] <= 16'b0100000011111110; //   SB R3, -2(R0)
      mem[27] <= 16'b0010010011000001; //   LB R3, 1(R2)
      mem[28] <= 16'b0100000011111111; //   SB R3, -1(R0)
      mem[29] <= 16'b0010000001111000; //   LB R1, -8(R0)
      mem[30] <= 16'b1111110000101000; //   ADD R5, R6, R0
      mem[31] <= 16'b1111111000110000; //   ADD R6, R7, R0
      mem[32] <= 16'b1111010000111000; //   ADD R7, R2, R0
      mem[33] <= 16'b1111110101001001; //   SUB R1, R6, R5
      mem[34] <= 16'b1111001000100000; //   ADD R4, R1, R0
      mem[35] <= 16'b1111111110001001; //   SUB R1, R7, R6
      mem[36] <= 16'b1111001000011000; //   ADD R3, R1, R0
      mem[37] <= 16'b1011100000000010; //   BLTZ R4, 2
      mem[38] <= 16'b1111100000101000; //   ADD R5, R4, R0
      mem[39] <= 16'b1000000000000010; //   BEQ R0, R0, 2
      mem[40] <= 16'b1111000100101001; //   SUB R5, R0, R4
      mem[41] <= 16'b1011011000000010; //   BLTZ R3, 2
      mem[42] <= 16'b1111011000110000; //   ADD R6, R3, R0
      mem[43] <= 16'b1000000000000010; //   BEQ R0, R0, 2
      mem[44] <= 16'b1111000011110001; //   SUB R6, R0, R3
      mem[45] <= 16'b1111101001001001; //   SUB R1, R5, R1
      mem[46] <= 16'b1011001000001010; //   BLTZ R1, 10
      mem[47] <= 16'b1111110001001001; //   SUB R1, R6, R1
      mem[48] <= 16'b1011001000001000; //   BLTZ R1, 8
      mem[49] <= 16'b1011100000000010; //   BLTZ R4, 2
      mem[50] <= 16'b1010011000000100; //   BGEZ R3, 4
      mem[51] <= 16'b1011011000000010; //   BLTZ R3, 2
      mem[52] <= 16'b1010100000000001; //   BGEZ R4, 1
      mem[53] <= 16'b1000000000000100; //   BEQ R0, R0, 4
      mem[54] <= 16'b0101000001011110; //   ADDI R1, R0, 30
      mem[55] <= 16'b0101001001001100; //   ADDI R1, R1, 12
      mem[56] <= 16'b1111001000001100; //   SLL R1, R1
      mem[57] <= 16'b1111001000001100; //   SLL R1, R1
      mem[58] <= 16'b0101001001000010; //   ADDI R1, R1, 2
      mem[59] <= 16'b0100000001111001; //   SB R1, -7(R0)
      mem[60] <= 16'b1000000000000010; //   BEQ R0, R0, 2
      mem[61] <= 16'b0101000001000000; //   ADDI R1, R0, 0
      mem[62] <= 16'b0100000001111001; //   SB R1, -7(R0)

      for(i = 63; i < 128; i = i + 1) begin
        mem[i] <= 16'b0000000000000000;
      end
    end
  end

endmodule
